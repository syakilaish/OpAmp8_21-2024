* Created by KLayout

* cell Op8_21
* pin Bias
* pin Out
* pin In-
* pin In+
* pin Vdd
* pin Vss
.SUBCKT Op8_21 1 7 10 12 14 24
* net 1 Bias
* net 7 Out
* net 10 In-
* net 12 In+
* net 14 Vdd
* net 24 Vss
* device instance $1 r0 *1 175,47.5 NMOS
M$1 7 6 24 24 NMOS L=1U W=96U AS=112P AD=112P PS=126U PD=126U
* device instance $7 m90 *1 95.5,41.5 NMOS
M$7 3 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $8 r0 *1 109.5,41.5 NMOS
M$8 4 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $9 m90 *1 47.5,41.5 NMOS
M$9 8 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $10 r0 *1 59,41.5 NMOS
M$10 2 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $11 r0 *1 124.5,40.5 NMOS
M$11 5 1 24 24 NMOS L=5U W=9U AS=16.5P AD=16.5P PS=23U PD=23U
* device instance $14 m90 *1 165.5,111.5 NMOS
M$14 18 15 6 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $19 m90 *1 164.5,49 NMOS
M$19 9 9 24 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $24 m90 *1 164.5,78 NMOS
M$24 15 15 9 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $29 m90 *1 95,61 NMOS
M$29 13 1 3 24 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $34 r0 *1 112,61 NMOS
M$34 6 1 4 24 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $39 r0 *1 55.5,56 NMOS
M$39 11 1 2 24 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $40 m90 *1 46,56 NMOS
M$40 1 1 8 24 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $41 m0 *1 180.5,95 PMOS
M$41 14 18 7 14 PMOS L=1U W=300U AS=420P AD=420P PS=434U PD=434U
* device instance $44 m90 *1 99.5,185.5 PMOS
M$44 22 19 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $49 r0 *1 113,185.5 PMOS
M$49 21 19 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $54 m90 *1 179,165.5 PMOS
M$54 17 17 14 14 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $61 r0 *1 79,104.5 PMOS
M$61 3 10 16 16 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $66 m90 *1 67.5,104.5 PMOS
M$66 4 12 16 16 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $71 r0 *1 156,183.5 PMOS
M$71 15 11 14 14 PMOS L=5U W=24U AS=48P AD=48P PS=52U PD=52U
* device instance $72 m90 *1 141.5,98.5 PMOS
M$72 6 5 18 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $82 m90 *1 154.5,149 PMOS
M$82 5 5 17 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $92 m90 *1 85,153.5 PMOS
M$92 19 13 22 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $97 r0 *1 96,153.5 PMOS
M$97 18 13 21 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $102 r0 *1 47.5,161 PMOS
M$102 16 11 23 14 PMOS L=2U W=40U AS=60P AD=60P PS=66U PD=66U
* device instance $104 r0 *1 49,188 PMOS
M$104 23 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $106 r0 *1 37.5,161 PMOS
M$106 11 11 20 14 PMOS L=2U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $107 m90 *1 36,188 PMOS
M$107 20 11 14 14 PMOS L=5U W=15U AS=30P AD=30P PS=34U PD=34U
* device instance $108 r0 *1 34.5,126.5 HRES
R$108 13 19 49000 HRES
* device instance $109 m0 *1 32,71 HRES
R$109 14 1 805000 HRES
* device instance $113 r0 *1 269.25,60 CAP
C$113 7 6 9.49e-13 CAP
* device instance $115 m0 *1 269.25,177.5 CAP
C$115 7 18 9.49e-13 CAP
.ENDS Op8_21
