* Created by KLayout

* cell Op8_21_V2_rev1
* pin Bias
* pin Out
* pin In-
* pin In+
* pin Vdd
* pin Vss
.SUBCKT Op8_21_V2_rev1 1 7 10 12 14 24
* net 1 Bias
* net 7 Out
* net 10 In-
* net 12 In+
* net 14 Vdd
* net 24 Vss
* device instance $1 r0 *1 175,47.5 NMOS
M$1 7 6 24 24 NMOS L=1U W=96U AS=112P AD=112P PS=126U PD=126U
* device instance $7 r0 *1 109.5,41.5 NMOS
M$7 4 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $8 m90 *1 95.5,41.5 NMOS
M$8 3 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $9 m90 *1 47.5,41.5 NMOS
M$9 8 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $10 r0 *1 59,41.5 NMOS
M$10 2 1 24 24 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $11 r0 *1 124.5,40.5 NMOS
M$11 5 1 24 24 NMOS L=5U W=9U AS=16.5P AD=16.5P PS=23U PD=23U
* device instance $14 m90 *1 95,61 NMOS
M$14 13 1 3 24 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $19 r0 *1 112,61 NMOS
M$19 6 1 4 24 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $24 r0 *1 55.5,56 NMOS
M$24 11 1 2 24 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $25 m90 *1 46,56 NMOS
M$25 1 1 8 24 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $26 m90 *1 165.5,111.5 NMOS
M$26 18 15 6 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $31 m90 *1 164.5,49 NMOS
M$31 9 9 24 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $36 m90 *1 164.5,78 NMOS
M$36 15 15 9 24 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $41 m90 *1 36,188 PMOS
M$41 21 11 14 14 PMOS L=5U W=15U AS=30P AD=30P PS=34U PD=34U
* device instance $42 r0 *1 37.5,161 PMOS
M$42 11 11 21 14 PMOS L=2U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $43 m0 *1 180.5,95 PMOS
M$43 14 18 7 14 PMOS L=1U W=300U AS=420P AD=420P PS=434U PD=434U
* device instance $46 m90 *1 99.5,185.5 PMOS
M$46 23 19 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $51 r0 *1 113,185.5 PMOS
M$51 20 19 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $56 m90 *1 179,165.5 PMOS
M$56 17 17 14 14 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $63 r0 *1 79,104.5 PMOS
M$63 3 10 16 16 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $68 m90 *1 67.5,104.5 PMOS
M$68 4 12 16 16 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $73 r0 *1 156,183.5 PMOS
M$73 15 11 14 14 PMOS L=5U W=24U AS=48P AD=48P PS=52U PD=52U
* device instance $74 m90 *1 141.5,98.5 PMOS
M$74 6 5 18 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $84 m90 *1 154.5,149 PMOS
M$84 5 5 17 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $94 m90 *1 85,153.5 PMOS
M$94 19 13 23 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $99 r0 *1 96,153.5 PMOS
M$99 18 13 20 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $104 r0 *1 47.5,161 PMOS
M$104 16 11 22 14 PMOS L=2U W=40U AS=60P AD=60P PS=66U PD=66U
* device instance $106 r0 *1 49,188 PMOS
M$106 22 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $108 r0 *1 21.05,135 HRES
R$108 13 19 50666.6666667 HRES
* device instance $109 m0 *1 35.65,73 HRES
R$109 1 14 800000 HRES
* device instance $117 r0 *1 274.25,60 CAP
C$117 7 6 1.022e-12 CAP
* device instance $119 m0 *1 274.25,177.5 CAP
C$119 7 18 1.022e-12 CAP
.ENDS Op8_21_V2_rev1
